library IEEE;
    use IEEE.std_logic_1164.all;
    use IEEE.numeric_std.all;

entity NewVhdlFile2 is
    port (
        clk: in  std_logic;
        rst: in  std_logic
    );
end entity;

architecture rtl of NewVhdlFile2 is
begin
end architecture;